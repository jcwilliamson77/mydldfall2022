module datapath2 ();

assign seed = ;

mux21 m1(seed, z_out, intial , y)

datapath d1(y, z)

flopr (z, z_out)

endmodule