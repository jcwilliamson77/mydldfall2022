module REG ();