module control_logic (clk, reset, seed, current_iteration, next_iteration);
    input logic [63:0] current_iteration;
    input logic clk;
    input logic reset;
    input logic [63:0] seed;
    output logic [63:0] next_iteration;
    logic [63:0] y;
    logic decision;


 
   
endmodule